`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:41:52 10/22/2019
// Design Name:   buffer_ram_dp
// Module Name:   C:/Users/UECCI/Documents/GitHub/SPARTAN6-ATMEGA-MAX5864/lab/P001-ProyectoCamara/src/ramdp/TB_ram.v
// Project Name:  P001-ProyectoCamara
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: buffer_ram_dp
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TB_ram;

	// Inputs
	reg clk;
	reg [16:0] addr_in;
	reg [15:0] data_in;
	reg regwrite;
	reg [16:0] addr_out;
	reg regread;

	// Outputs
	wire [15:0] data_out;
	
	//Simulation registers
	reg [4:0] DR;
	reg [5:0] DG;
	reg [4:0] DB;

	// Instantiate the Unit Under Test (UUT)
	buffer_ram_dp uut (
		.clk(clk), 
		.addr_in(addr_in), 
		.data_in(data_in), 
		.regwrite(regwrite), 
		.data_out(data_out), 
		.addr_out(addr_out), 
		.regread(regread)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		addr_in = 0;
		data_in = 0;
		regwrite = 0;
		addr_out = 0;
		regread = 1;
		
		DR=0;
		DG=0;
		DB=0;

  // Adicionar las estimulos necesarios para simular la lectura y escritura de la memoria ram
		for(addr_out=0; addr_out<65535; addr_out=addr_out+1) begin
			//Nueva Addrress
			addr_in = addr_out;
			#2;//Espera a lectura
			regread = 0;
			//Ingrese nuevo codigo de Color
			DG=DG+8;
			if(DG==0)begin
				DR=DR+4;
				if(DR==0)
					DB=DB+4;
			end
			data_in = {DR,DG,DB};
			regwrite = 1;
			#2;//Espera a escritura
			regwrite = 0;
			regread = 1;
			#2;//Espera a segunda lectura
		end
		
	end
	
	always #1 clk = ~clk ;
	
endmodule

